//===================================================================================
// Project      : aes (advanced encryption standard)
// File name    : key_exp_top.sv 
// Designer     : Albin Gomes
// Device       : 
// Description  :
// Limitations  :
// Version      :
//===================================================================================

module key_exp_top (
  // Input
  input           clk,
  input           reset_n,
  input [4:0]     round,
  input [127:0]   key,
  // Output
  output[127:0]  key_out
);

//-----------------------------------------------------------------------------------
// Nets and Regs
//-----------------------------------------------------------------------------------




















endmodule