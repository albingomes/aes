//===================================================================================
// Project      : aes (advanced encryption standard)
// File name    : g_function.sv 
// Designer     : Albin Gomes
// Device       : 
// Description  :
// Limitations  :
// Version      :
//===================================================================================

module g_function (
  input           clk,
  input           reset_n,
  input           enable,
  input   [31:0]  data_in,
  output  [31:0]  data_out,
  output          done
);






endmodule