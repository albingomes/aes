//===================================================================================
// Project      : aes (advanced encryption standard)
// File name    : s_box.sv 
// Designer     : Albin Gomes
// Device       : 
// Description  :
// Limitations  :
// Version      :
//===================================================================================

module s_box (
  input         clk,
  input         reset_n,
  input         enable,
  input   [7:0] data_in,
  output  [7:0] data_out,
  output        done
);

//-----------------------------------------------------------------------------------
// Nets, Regs and states
//-----------------------------------------------------------------------------------

//-----------------------------------------------------------------------------------
// Instantiations
//-----------------------------------------------------------------------------------

//-----------------------------------------------------------------------------------
// Assignment
//-----------------------------------------------------------------------------------

//-----------------------------------------------------------------------------------
// Process
//-----------------------------------------------------------------------------------



endmodule